VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.001 ;

PROPERTYDEFINITIONS
LAYER LEF58_NOCUTCLASS STRING ;
LAYER LEF58_AREA STRING ;
LAYER LEF58_ARRAYSPACING STRING ;
LAYER LEF58_BOUNDARYBLOCKAGE STRING ;
LAYER LEF58_BOUNDARYEOLBLOCKAGE STRING ;
LAYER LEF58_COREEOLBLOCKAGE STRING ;
LAYER LEF58_CORNEREOLKEEPOUT STRING ;
LAYER LEF58_CORNERFILLSPACING STRING ;
LAYER LEF58_CORNERSPACING STRING ;
LAYER LEF58_CUTCLASS STRING ;
LAYER LEF58_CUTONCENTERLINE STRING ;
LAYER LEF58_ENCLOSUREEDGE STRING ;
LAYER LEF58_ENCLOSURESPACING STRING ;
LAYER LEF58_ENCLOSURE STRING ;
LAYER LEF58_KEEPOUTZONE STRING ;
LAYER LEF58_DIRECTIONALSPACING STRING ;
LAYER LEF58_ENCLOSURETABLE STRING ;
LAYER LEF58_ENCLOSURETOJOINT STRING ;
LAYER LEF58_ENCLOSUREWIDTH STRING ;
LAYER LEF58_ENCLOSUREWITHEOL STRING ;
LAYER LEF58_EOLENCLOSURE STRING ;
LAYER LEF58_EOLEXTENSIONSPACING STRING ;
LAYER LEF58_EOLKEEPOUT STRING ;
LAYER LEF58_EOLTRACK STRING ;
LAYER LEF58_FILLTOFILLSPACING STRING ;
LAYER LEF58_FIVEWIRESEOLSPACING STRING ;
LAYER LEF58_FORBIDDENSPACING STRING ;
LAYER LEF58_GAP STRING ;
LAYER LEF58_JOINTCORNERSPACING STRING ;
LAYER LEF58_LINEENDGAP STRING ;
LAYER LEF58_LITHOMACROHALO STRING ;
LAYER LEF58_MAXSPACING STRING ;
LAYER LEF58_MAXWIDTH STRING ;
LAYER LEF58_MINIMUMCUT STRING ;
LAYER LEF58_MINLENGTHPARALLEL STRING ;
LAYER LEF58_MINSIZE STRING ;
LAYER LEF58_MINSTEP STRING ;
LAYER LEF58_OPPOSITEEOLSPACING STRING ;
LAYER LEF58_OPPOSITEOVERLAPCUTSPACING STRING ;
LAYER LEF58_PINCONNECTBLOCKAGE STRING ;
LAYER LEF58_PITCH STRING ;
LAYER LEF58_PROTRUSIONWIDTH STRING ;
LAYER LEF58_RECTONLY STRING ;
LAYER LEF58_REGION STRING ;
LAYER LEF58_RIGHTWAYONGRIDONLY STRING ;
LAYER LEF58_SAMEMETALALIGNEDCUTS STRING ;
LAYER LEF58_SPACING STRING ;
LAYER LEF58_SPACINGTABLE STRING ;
LAYER LEF58_SPANLENGTHENCLOSURESPACING STRING ;
LAYER LEF58_SPANLENGTHTABLE STRING ;
LAYER LEF58_TWOWIRESFORBIDDENSPACING STRING ;
LAYER LEF58_TYPE STRING ;
LAYER LEF58_VOLTAGESPACING STRING ;
LAYER LEF58_WIDTHTABLE STRING ;
LAYER LEF58_WRNGDIREOLKEEPOUT STRING ;
END PROPERTYDEFINITIONS

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER Gate
  TYPE MASTERSLICE ;
END Gate

LAYER Active
  TYPE MASTERSLICE ;

END Active

LAYER V0
  TYPE CUT ;
  SPACING 0.072 ;
  WIDTH 0.072 ;
END V0

LAYER M1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.144 ;
  WIDTH 0.072 ;
  SPACING 0.072 ;
  AREA 0.010656 ;                   # Min Area # This should ideally be 16x not 4x as each dimension is scaled up by 16
                                    # we only allow landing on pins (set in router) so area should not matter
  SPACING 0.072 RANGE 0.144 4.000 ; # This rule is redundant with the SPACING rule

  PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.073 EXTENSION 0 0 0.124 ;" ; #  Tip to Tip Spacing
OFFSET 0.0 ;
  PROPERTY LEF58_CORNERSPACING "CORNERSPACING CONVEXCORNER CORNERONLY 0.040 WIDTH 0.072 SPACING 0.072 ;" ;
PROPERTY LEF58_AREA "AREA 0.017 EXCEPTSTEP 0.12 0.05 ; " ;
PROPERTY LEF58_BOUNDARYBLOCKAGE " BOUNDARYBLOCKAGE 0.02 ; " ;
PROPERTY LEF58_MAXWIDTH " MAXWIDTH  0.12 ; " ;
PROPERTY LEF58_CORNERSPACING  " CORNERSPACING CONVEXCORNER CORNERONLY 0.050 WIDTH 0.000 SPACING 0.100 ; " ;
PROPERTY LEF58_EOLEXTENSIONSPACING "EOLEXTENSIONSPACING 0.1 ENDOFLINE 0.11 EXTENSION 0.14 ENDOFLINE 0.15 EXTENSION 0.12 ENDTOEND 0.13 ; " ;
PROPERTY LEF58_EOLKEEPOUT "EOLKEEPOUT 0.2 EXTENSION 0.03 0.05 0.1 ; " ;
PROPERTY LEF58_FORBIDDENSPACING "FORBIDDENSPACING 0.01 0.25 WIDTH 0.05 PRL 0.15 ; " ;
PROPERTY LEF58_GAP " GAP EXACTWIDTH 0.2 MAXLENGTH 0.6 SPACING 0 0.4 1 0.3 2 0.5 ENDTOEND 0.8 ; " ;
PROPERTY LEF58_JOINTCORNERSPACING "JOINTCORNERSPACING 0.05 JOINTWIDTH 0.07 JOINTLENGTH 0.06 EDGELENGTH 0.1 ; " ;
PROPERTY LEF58_MINIMUMCUT "MINIMUMCUT 2 WIDTH 0.2 SAMEMETALOVERLAP ; " ;
PROPERTY LEF58_MINSTEP "MINSTEP 0.5 MAXEDGES 1 NOBETWEENEOL 1.0 ; " ;
PROPERTY LEF58_PITCH " PITCH 0.1 FIRSTLASTPITCH 0.14 ; " ;
PROPERTY LEF58_PROTRUSIONWIDTH "PROTRUSIONWIDTH 0.05 WIDTH 0.11 MINLENGTH 0.12 WIDTH 0.15 MINLENGTH 0.14 ; " ;  
PROPERTY LEF58_RECTONLY   " RECTONLY ; " ;
PROPERTY LEF58_SPANLENGTHTABLE   " SPANLENGTHTABLE 0.05 0.06 0.07 0.080 0.090 0.10 ; SPANLENGTHTABLE 0.07 0.10 WRONGDIRECTION EXCEPTOTHERSPAN 0.05 ; " ;
PROPERTY LEF58_SPACING "SPACING 0.15 AREA 0.03 ; " ;
PROPERTY LEF58_TWOWIRESFORBIDDENSPACING  " TWOWIRESFORBIDDENSPACING SAMEMASK 0.02 0.20 MINSPANLENGTH 0.05 EXACTSPANLENGTH MAXSPANLENGTH 0.08 EXACTSPANLENGTH PRL 0 ; " ;
END M1

LAYER V1
  TYPE CUT ;
  SPACING 0.072 ;     # unlike generate, this is really spacing, not center to center.
  WIDTH 0.072 ;
PROPERTY LEF58_ARRAYSPACING  " ARRAYSPACING WITHIN 0.2 ARRAYWIDTH 0.06 CUTSPACING 0.05 ARRAYCUTS 3 SPACING 0.05 ; " ;
PROPERTY LEF58_ENCLOSURE " ENCLOSURE  0.03 0.03 WIDTH 0.3 EXCEPTEXTRACUT 0.2 ; " ;
PROPERTY LEF58_ENCLOSUREEDGE "ENCLOSUREEDGE 0.02 WIDTH 0.2 PARALLEL 0.25 WITHIN 0.11 ; " ;
PROPERTY LEF58_ENCLOSURETABLE "ENCLOSURETABLE WIDTH 0.3 0.05 0.05 0.08 0.1; " ;
PROPERTY LEF58_ENCLOSURETOJOINT "ENCLOSURETOJOINT 0.05 0.03 JOINTWIDTH 0.15 JOINTLENGTH 0.1 ; " ;
PROPERTY LEF58_SPACING "SPACING 0.15 SAMEMASK ; " ;
PROPERTY LEF58_ENCLOSUREEDGE "ENCLOSUREEDGE ABOVE 0.02 OPPOSITE ; " ;
PROPERTY LEF58_OPPOSITEOVERLAPCUTSPACING " OPPOSITEOVERLAPCUTSPACING 0.06 PRL 0.01 LAYER M1 ; " ;
END V1

LAYER M2
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  WIDTH 0.072 ; # Min Width
  SPACING 0.072 ; # Min Spacing

  OFFSET -1.080 ;

  #  MINSIZE is set so that the minimum lenght of a segment is 36nm. At the proper rule size of
  #  31nm, the lines can't be minimum space. This causes DRCs (like crazy). Same for M3
  #  MINSIZE 0.112 0.072 ;
  # area is adjusted to match this (Nanoroute requires both AREA and MINSIZE)

  AREA 0.010656 ;
  MINSIZE 0.148 0.072 ;

  PITCH 0.180 0.144 ;

  # this enforces the correct routing tracks on M2 with wide M2 power rails

  PROPERTY LEF58_PITCH "
   PITCH 0.144 FIRSTLASTPITCH 0.180
   ;
  " ;

  # this checks for distance in any direction so is not correct
  # 0.070 is to avoid conflicts with the adjacent lines. This should be caught by CORNERSPACING below
  #   SPACING 0.124 ENDOFLINE 0.1 WITHIN 0.070 ;

  PROPERTY LEF58_SPACING
    " SPACING 0.072 ENDOFLINE 0.1 WITHIN 0.08 ENDTOEND 0.124
      PARALLELEDGE 0.100 WITHIN 0.08 ; " ;  

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.0 0.05 0.124 CORNERONLY ;
  " ;

  PROPERTY LEF58_CORNERSPACING "
     CORNERSPACING CONVEXCORNER WIDTH 0.000 SPACING 0.080 ;
  " ; # CORNER to CORNER SPACING Rule

  # Originally no width table for M2 since it is the follow rails.
  # They can be 1x or 2x (2x causes DRCs on SAV V1). However, this seems to allow a double width M2
  # on vias, which violates. Thus, this is added. Note that wide power follow rails will violate.

  PROPERTY LEF58_WIDTHTABLE "
      WIDTHTABLE 0.072 0.36 0.648 0.936 1.224 1.512 ;
  " ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;
  PROPERTY LEF58_CORNEREOLKEEPOUT
     " CORNEREOLKEEPOUT WIDTH 0.1
          EOLSPACING 0.124
          EXTENSION 0.08 0.094 0.08 ; " ;

END M2

LAYER V2
  TYPE CUT ;
  SPACING 0.072 ;
  WIDTH 0.072 ;

  # V1.LW.1, V1PWR.LW.1, V1BAR.LW.1, V1LRG.LW.1
  PROPERTY LEF58_CUTCLASS "
    CUTCLASS Vx    WIDTH 0.020 LENGTH 0.020 CUTS 1 ;
    CUTCLASS VxPWR WIDTH 0.020 LENGTH 0.030 CUTS 1 ;
    CUTCLASS VxBAR WIDTH 0.020 LENGTH 0.040 CUTS 2 ;
    CUTCLASS VxLRG WIDTH 0.040 LENGTH 0.040 CUTS 4 ; " ;

  # V1.S.2
  PROPERTY LEF58_MAXSPACING "
    MAXSPACING 1.000 CUTCLASS Vx ; " ;

  # V1.S.1/5, V1PWR.S.V1.1, V1.S.V1BAR.1, V1.S.V1LRG.1
  # V1PWR.S.1, V1PWR.S.V1BAR.1, V1PWR.S.V1LRG.1/2
  # V1BAR.S.1/2/3, V1BAR.S.V1LRG.1/2  
  # V1LRG.S.1  
  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
    CENTERTOCENTER Vx TO Vx  Vx TO VxLRG  VxLRG TO VxLRG
    CENTERANDEDGE VxBAR TO VxLRG VxPWR TO VxLRG
    EXACTALIGNEDSPACING Vx 0.034      
    CUTCLASS        Vx               VxPWR SIDE     VxPWR END      VxBAR SIDE     VxBAR END      VxLRG
    Vx            0.045    0.045   0.02475 0.042  0.02475 0.042  0.0415 0.0415  0.0415 0.0415  0.130 0.130
    VxPWR SIDE    0.02475  0.042   0.042 0.042    0.042 0.042    0.042 0.042    0.042 0.042    0.100 0.130
    VxPWR END     0.02475  0.042   0.042 0.042    0.042 0.042    0.042 0.042    0.042 0.042    0.124 0.130
    VxBAR SIDE    0.0415   0.0415  0.042 0.042    0.042 0.042    0.042 0.042    0.042 0.042    0.100 0.130
    VxBAR END     0.0415   0.0415  0.042 0.042    0.042 0.042    0.042 0.042    0.042 0.042    0.124 0.130
    VxLRG         0.130    0.130   0.100 0.130    0.124 0.130    0.100 0.130    0.124 0.130    0.160 0.160 ; " ;

PROPERTY LEF58_CUTCLASS "CUTCLASS Vx WIDTH 0.15 ; " ;  
PROPERTY LEF58_FORBIDDENSPACING "FORBIDDENSPACING CUTCLASS Vx 0.07 0.09 SHORTEDGEONLY ; " ;
PROPERTY LEF58_NOCUTCLASS "NOCUTCLASS Vx EXCEPTMULTICUTS ; " ;
PROPERTY LEF58_SAMEMETALALIGNEDCUTS "SAMEMETALALIGNEDCUTS 2 CUTCLASS ALL BELOW WIDTH 0.04 SPACING 0.1 ; " ;

END V2

LAYER M3
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.144 ;
  OFFSET 0.0 ;
  WIDTH 0.072 ; # Min Width
  SPACING 0.072 ; # Min Spacing

  #  MINSIZE is set so that the minimum lenght of a segment is 36nm. At the proper rule size of
  #  31nm, the lines can't be minimum space. This causes DRCs (like crazy). Same for M2
  #  MINSIZE 0.112 0.072 ;
  # area is adjusted to match this (Nanoroute requires both AREA and MINSIZE)

  AREA 0.010656 ;
  MINSIZE 0.148 0.072 ;

  PROPERTY LEF58_SPACING
    " SPACING 0.072 ENDOFLINE 0.1 WITHIN 0.05 ENDTOEND 0.124  
      PARALLELEDGE 0.100 WITHIN 0.08 ; " ;  

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.0 0.05 0.124 CORNERONLY ;
  " ;

  PROPERTY LEF58_CORNERSPACING "
   CORNERSPACING CONVEXCORNER WIDTH 0.000 SPACING 0.080
   ;
  " ; # CORNER to CORNER SPACING Rule

  # to make the special route widths integer values of the tracks, i.e., 1, 5, 9, 13... min widths
  # the widths should be calculated in the APR tool, since viaGen does not seem to respect these

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.072 0.36 0.648 0.936 1.224 1.512 ; " ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M3

LAYER V3
  TYPE CUT ;

  # different format to allow long vias for SAV power connections

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS V3       WIDTH 0.072 LENGTH 0.096 CUTS 1  ;
    CUTCLASS V3_0p480 WIDTH 0.072 LENGTH 0.480 CUTS 4  ;
    CUTCLASS V3_0p864 WIDTH 0.072 LENGTH 0.864 CUTS 8  ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   V3 V3_0p480 V3_0p864
        V3       -  -        -        -  - -
        V3_0p480 -  -        -        -  - -
        V3_0p864 -  -        -        -  - -
    ;
  " ;

  # covered below?
  # ENCLOSURE CUTCLASS V3       END 0.02 SIDE 0.0 ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS V3 BELOW EOL 0.0 0.020 0.0 ;
    ENCLOSURE CUTCLASS V3 ABOVE EOL 0.0 0.044 0.0 ;
    ENCLOSURE CUTCLASS V3_0p480 END 0.0  SIDE 0.0 ;
    ENCLOSURE CUTCLASS V3_0p864 END 0.0  SIDE 0.0 ;
  " ;

  PROPERTY LEF58_KEEPOUTZONE "
     KEEPOUTZONE CUTCLASS V3 TO V3
        EXCEPTEXACTALIGNED 0.072
        HORIZONTALEXTENSION 0.092 0.092
        VERTICALEXTENSION 0.102 0.102
        SPIRALEXTENSION 0.112
  ; " ;
  PROPERTY LEF58_DIRECTIONALSPACING "
     DIRECTIONALSPACING 0.071 VERTICAL PRL 0.072
     CUTCLASS V3 TO V3 PARALLEL 0.071 WITHIN 0.072
  ; " ;

PROPERTY LEF58_ARRAYSPACING  " ARRAYSPACING WITHIN 0.2 ARRAYWIDTH 0.06 CUTSPACING 0.05 ARRAYCUTS 3 SPACING 0.05 ; " ;
PROPERTY LEF58_CUTONCENTERLINE "CUTONCENTERLINE 0.13 CUTCLASS V3 ; " ;
PROPERTY LEF58_ENCLOSURE " ENCLOSURE CUTCLASS V3 0.10 0.10 ; " ;
PROPERTY LEF58_MAXSPACING "MAXSPACING 0.01 CUTCLASS V3 ; " ;
PROPERTY LEF58_SPACING "SPACING 0.15 SAMEMASK ; " ;
PROPERTY LEF58_OPPOSITEOVERLAPCUTSPACING " OPPOSITEOVERLAPCUTSPACING 0.06 PRL 0.01 LAYER M1 ; " ;
PROPERTY LEF58_SAMEMETALALIGNEDCUTS "SAMEMETALALIGNEDCUTS 1 CUTCLASS ALL BELOW WIDTH 0.04 SPACING 0.1 ; " ;

END V3

LAYER M4
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.192 ;
  WIDTH 0.096 ;
  SPACING 0.096 ;

  OFFSET 0.012 ;

  AREA 0.032 ;

  PROPERTY LEF58_SPACING "
    SPACING 0.096 ENDOFLINE 0.1 WITHIN 0.160 ENDTOEND 0.160 ; " ;  

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.096 0.480 0.864 1.248 1.632 ; " ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.192
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.192 0.097 0.192 CORNERONLY ;
  " ;

  # spacing table is required for the rule that has wide metal requires a 72nm (288 scaled)
  # spacing between wide and minimum metals

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M4

LAYER V4
  TYPE CUT ;

  # spacing is 4 * 34 = 136
  # SPACING 0.136 ;
  # WIDTH 0.072 ;
  # ENCLOSURE 0.044 0.0 ;

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS Vx       WIDTH 0.096 LENGTH 0.096 ;
    CUTCLASS Vx_0p480 WIDTH 0.096 LENGTH 0.480 CUTS 4  ;
    CUTCLASS Vx_0p864 WIDTH 0.096 LENGTH 0.864 CUTS 8  ;
    CUTCLASS Vx_1p248 WIDTH 0.096 LENGTH 1.248 CUTS 12 ;
    CUTCLASS Vx_1p632 WIDTH 0.096 LENGTH 1.632 CUTS 16 ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
        Vx       -  -        -        -        - -  -        -        -        -
        Vx_0p480 -  -        -        -        - -  -        -        -        -
Vx_0p864 -  -        -        -        - -  -        -        -        -
Vx_1p248 -  -        -        -        - -  -        -        -        -
Vx_1p632 -  -        -        -        - -  -        -        -        -
    ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS Vx 0.044 0.0 ;
    ENCLOSURE CUTCLASS Vx EOL   0.0 0.044 0.044 ;
    ENCLOSURE CUTCLASS Vx_0p480 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_0p864 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p248 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p632 END 0.00 SIDE 0.0 ;
  " ;

END V4

LAYER M5
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.192 ;
  WIDTH 0.096 ;
  SPACING 0.096 ;
  OFFSET 0.0 ;

  AREA 0.032 ;

  PROPERTY LEF58_SPACING "
    SPACING 0.096 ENDOFLINE 0.1 WITHIN 0.160 ENDTOEND 0.160 ; " ;  

  MINIMUMDENSITY 60 ;
  MAXIMUMDENSITY 360 ;
  DENSITYCHECKWINDOW 80 80 ;
  DENSITYCHECKSTEP 40 ;

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.096 0.480 0.864 1.248 1.632 2.016 2.400 2.784 3.168 3.552 3.936 ; " ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.192
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.1 EXTENSION 0.192 0.097 0.192
    CORNERONLY ;
  " ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M5

LAYER V5
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS Vx       WIDTH 0.096 LENGTH 0.128 ;
    CUTCLASS Vx_0p480 WIDTH 0.096 LENGTH 0.640 CUTS 4  ;
    CUTCLASS Vx_0p864 WIDTH 0.096 LENGTH 1.152 CUTS 8  ;
    CUTCLASS Vx_1p248 WIDTH 0.096 LENGTH 1.664 CUTS 12 ;
    CUTCLASS Vx_1p632 WIDTH 0.096 LENGTH 2.176 CUTS 16 ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   Vx Vx_0p480 Vx_0p864 Vx_1p248 Vx_1p632
        Vx       -  -        -        -        - -  -        -        -        -
        Vx_0p480 -  -        -        -        - -  -        -        -        -
Vx_0p864 -  -        -        -        - -  -        -        -        -
Vx_1p248 -  -        -        -        - -  -        -        -        -
Vx_1p632 -  -        -        -        - -  -        -        -        -
    ;
  " ;

  # end refers to the end of the VIA! Thus, since it is rectangular the proper
  # enclosure is on the side not the end...
  # ENCLOSURE CUTCLASS Vx END 0.0 SIDE 0.044 ;  But--this refers to top and bottom
  # actually passing the rule is done by having the correct vias below.

  PROPERTY LEF58_ENCLOSURE "
  ENCLOSURE CUTCLASS Vx EOL 0.0 0.044 0.044 ;
  ENCLOSURE CUTCLASS Vx_0p480 END 0.00 SIDE 0.0 ;
  ENCLOSURE CUTCLASS Vx_0p864 END 0.00 SIDE 0.0 ;
  ENCLOSURE CUTCLASS Vx_1p248 END 0.00 SIDE 0.0 ;
  ENCLOSURE CUTCLASS Vx_1p632 END 0.00 SIDE 0.0 ;
  " ;


END V5

LAYER M6
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.256 ;
  WIDTH 0.128 ;
  SPACING 0.128 ;

  AREA 0.035 ;   # Areas still need tweaking

  PROPERTY LEF58_SPACING
    " SPACING 0.128 ENDOFLINE 0.15 WITHIN 0.160 ENDTOEND 0.160 ; " ;  

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.128 0.640 1.152 1.664 2.176 ; " ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.192
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.2 EXTENSION 0.192 0.129 0.192 CORNERONLY ;
  " ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M6

LAYER V6
  TYPE CUT ;

  PROPERTY LEF58_CUTCLASS "  
    CUTCLASS Vx       WIDTH 0.128 LENGTH 0.128 ;
    CUTCLASS Vx_0p640 WIDTH 0.128 LENGTH 0.640 CUTS 4  ;
    CUTCLASS Vx_1p152 WIDTH 0.128 LENGTH 1.152 CUTS 8  ;
    CUTCLASS Vx_1p664 WIDTH 0.128 LENGTH 1.664 CUTS 12 ;
    CUTCLASS Vx_2p176 WIDTH 0.128 LENGTH 2.176 CUTS 16 ;
  " ;

  PROPERTY LEF58_SPACINGTABLE "
    SPACINGTABLE
      DEFAULT 0.136
      CUTCLASS   Vx Vx_0p640 Vx_1p152 Vx_1p664 Vx_2p176
        Vx       -  -        -        -        - -  -        -        -        -
        Vx_0p640 -  -        -        -        - -  -        -        -        -
Vx_1p152 -  -        -        -        - -  -        -        -        -
Vx_1p664 -  -        -        -        - -  -        -        -        -
Vx_2p176 -  -        -        -        - -  -        -        -        -
    ;
  " ;

  PROPERTY LEF58_ENCLOSURE "
    ENCLOSURE CUTCLASS Vx 0.044  0.0 ;
    ENCLOSURE CUTCLASS Vx EOL 0.0 0.044 0.044 ;
    ENCLOSURE CUTCLASS Vx_0p640 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p152 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_1p664 END 0.00 SIDE 0.0 ;
    ENCLOSURE CUTCLASS Vx_2p176 END 0.00 SIDE 0.0 ;
  " ;

END V6

LAYER M7
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.256 ;
  WIDTH 0.128 ;
  SPACING 0.128 ;

  AREA 0.035 ;   # Areas still need tweaking

  PROPERTY LEF58_SPACING
    " SPACING 0.120 ENDOFLINE 0.15 WITHIN 0.160 ENDTOEND 0.160 ; " ;  

  PROPERTY LEF58_WIDTHTABLE
      " WIDTHTABLE 0.128 0.640 1.152 1.664 2.176 ; " ;
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PROPERTY LEF58_CORNERSPACING "
    CORNERSPACING CONVEXCORNER CORNERONLY 0.300
      WIDTH 0.000 SPACING 0.160 ;
  " ;

  PROPERTY LEF58_EOLKEEPOUT "
    EOLKEEPOUT 0.2 EXTENSION 0.192 0.129 0.192
    CORNERONLY ;
  " ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0.00
      WIDTH 0.000     0.096
      WIDTH 0.100     0.288 ;

  PROPERTY LEF58_RIGHTWAYONGRIDONLY "
      RIGHTWAYONGRIDONLY ;
  " ;

  PROPERTY LEF58_RECTONLY "
      RECTONLY ;
  " ;

END M7

LAYER V7
  TYPE CUT ;
  SPACING 0.184 ;
  WIDTH 0.128 ;
END V7

LAYER M8
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.32 0.32 ;
  WIDTH 0.16 ;
  AREA 30.08 ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.599 4.799 7.199
    WIDTH 0 0.16 0.16 0.16 0.16
    WIDTH 0.239 0.16 0.16 0.16 0.16
    WIDTH 0.319 0.16 0.16 0.16 0.16
    WIDTH 0.479 0.16 0.16 0.16 0.16
    WIDTH 1.999 0.16 0.16 0.16 2
    WIDTH 3.999 0.16 0.16 0.16 4 ;

  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMABOVE ;
  MAXWIDTH 8 ;
  MINSTEP 0.16 STEP ;
END M8

LAYER V8
  TYPE CUT ;
  SPACING 0.228 ;
  WIDTH 0.16 ;
END V8


LAYER M9
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.32 0.32 ;
  WIDTH 0.16 ;
  AREA 30.08 ;

  SPACINGTABLE
    PARALLELRUNLENGTH 0 1.599 4.799 7.199
    WIDTH 0 0.16 0.16 0.16 0.16
    WIDTH 0.239 0.16 0.16 0.16 0.16
    WIDTH 0.319 0.16 0.16 0.16 0.16
    WIDTH 0.479 0.16 0.16 0.16 0.16
    WIDTH 1.999 0.16 0.16 0.16 2
    WIDTH 3.999 0.16 0.16 0.16 4 ;

  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMABOVE ;
  MINSTEP 0.16 STEP ;
END M9

LAYER V9
  TYPE CUT ;
  SPACING 0.228 ;
  WIDTH 0.16 ;
END V9

LAYER Pad
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.32 0.32 ;
  WIDTH 0.16 ;
  SPACINGTABLE
    PARALLELRUNLENGTH 0 47.999
    WIDTH 0 8 8
    WIDTH 47.999 8 12 ;
  MINIMUMCUT 1 WIDTH 0.16 WITHIN 6.82 FROMBELOW ;
  MINIMUMCUT 1 WIDTH 1.44 WITHIN 6.82 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 7.22 WITHIN 6.82 FROMBELOW ;
  MINIMUMDENSITY 80 ;
  MAXIMUMDENSITY 320 ;
  DENSITYCHECKWINDOW 400 400 ;
  DENSITYCHECKSTEP 200 ;
END Pad


VIA VIA9Pad Default
  LAYER M9 ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER Pad ;
    RECT -0.2 -0.2 0.2 0.2 ;
  LAYER V9 ;
    RECT -0.2 -0.2 0.2 0.2 ;
END VIA9Pad

VIA VIA89 Default
  LAYER M8 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER M9 ;
    RECT -0.08 -0.08 0.08 0.08 ;
  LAYER V8 ;
    RECT -0.08 -0.08 0.08 0.08 ;
END VIA89

VIA VIA78 Default
  LAYER M7 ;
    RECT -0.064 -0.108 0.064 0.108 ;
  LAYER M8 ;
    RECT -0.108 -0.080 0.108 0.080 ;
  LAYER V7 ;
    RECT -0.064 -0.064 0.064 0.064 ;
END VIA78

VIA VIA67 Default
  LAYER M6 ;
    RECT -0.108 -0.064 0.108 0.064 ;
  LAYER M7 ;
    RECT -0.064 -0.108 0.064 0.108 ;
  LAYER V6 ;
    RECT -0.064 -0.064 0.064 0.064 ;
END VIA67

VIA VIA56 Default
  LAYER M5 ;
    RECT -0.048 -0.108 0.048 0.108 ;
  LAYER M6 ;
    RECT -0.092 -0.064 0.092 0.064 ;
  LAYER V5 ;
    RECT -0.048 -0.064 0.048 0.064 ;
END VIA56

VIA VIA45 Default
  LAYER M4 ;
    RECT -0.092 -0.048 0.092 0.048 ;
  LAYER M5 ;
    RECT -0.048 -0.092 0.048 0.092 ;
  LAYER V4 ;
    RECT -0.048 -0.048 0.048 0.048 ;
END VIA45

VIA VIA34 Default
  LAYER M3 ;
    RECT -0.036 -0.068 0.036 0.068 ;
  LAYER M4 ;
    RECT -0.080 -0.048 0.080 0.048 ;
  LAYER V3 ;
    RECT -0.036 -0.048 0.036 0.048 ;
END VIA34

VIA VIA23 Default
  LAYER M2 ;
    RECT -0.056 -0.036 0.056 0.036 ;
  LAYER M3 ;
    RECT -0.036 -0.056 0.036 0.056 ;
  LAYER V2 ;
    RECT -0.036 -0.036 0.036 0.036 ;
END VIA23

VIA VIA12 Default
  LAYER M1 ;
    RECT -0.036 -0.044 0.036 0.044 ;
  LAYER M2 ;
    RECT -0.056 -0.036 0.056 0.036 ;
  LAYER V1 ;
    RECT -0.036 -0.036 0.036 0.036 ;
END VIA12


END LIBRARY
